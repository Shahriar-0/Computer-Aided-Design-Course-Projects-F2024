module DP(input clk, rst, ld1, ld2, ld3, ld4);

    

endmodule