module AND2 (
    input A, B,

    output out
);

    __ACT_C1 and3(0, 0, 0, 0, 1, B, A, 0, out);

endmodule