module NOT (
    input A,
    
    output out
);

    __ACT_C1 not(1, 1, 1, 0, 0, 0, 0, A, out);

endmodule