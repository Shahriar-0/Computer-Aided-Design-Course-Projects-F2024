module AND4 (
    input A0, A1, B0, B1,

    output out
);

    __ACT_C2 and4(0, 0, 0, A1, 0, B1, A0, B0, out); 

endmodule