module AND3 (
    input A, B, C,

    output out
);

    __ACT_C1 and3(0, 0, 0, 0, A, B, C, 0, out);

endmodule